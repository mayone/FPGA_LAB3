module circle(center_x, center_y, R, G, B,);

        input center;
        
endmodule
