module circle(center);

        input center;
        
endmodule
