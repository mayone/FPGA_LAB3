module circle(center_x, center_y, HSYNC, VSYNC, R, G, B);

        input   center_x, center_y;
        output  HSYNC, VSYNC;
        output  R, G, B;

        // variables
        
        // design
        
endmodule
